netcdf \20210305T1600Z-B20210303T0600Z-temperature_at_screen_level {
dimensions:
	threshold = 63 ;
	projection_y_coordinate = 970 ;
	projection_x_coordinate = 1042 ;
	bnds = 2 ;
variables:
	float probability_of_air_temperature_above_threshold(threshold, projection_y_coordinate, projection_x_coordinate) ;
		probability_of_air_temperature_above_threshold:least_significant_digit = 3LL ;
		probability_of_air_temperature_above_threshold:long_name = "probability_of_air_temperature_above_threshold" ;
		probability_of_air_temperature_above_threshold:units = "1" ;
		probability_of_air_temperature_above_threshold:grid_mapping = "lambert_azimuthal_equal_area" ;
		probability_of_air_temperature_above_threshold:coordinates = "blend_time forecast_period forecast_reference_time height time" ;
	int lambert_azimuthal_equal_area ;
		lambert_azimuthal_equal_area:grid_mapping_name = "lambert_azimuthal_equal_area" ;
		lambert_azimuthal_equal_area:longitude_of_prime_meridian = 0. ;
		lambert_azimuthal_equal_area:semi_major_axis = 6378137. ;
		lambert_azimuthal_equal_area:semi_minor_axis = 6356752.31414036 ;
		lambert_azimuthal_equal_area:longitude_of_projection_origin = -2.5 ;
		lambert_azimuthal_equal_area:latitude_of_projection_origin = 54.9 ;
		lambert_azimuthal_equal_area:false_easting = 0. ;
		lambert_azimuthal_equal_area:false_northing = 0. ;
	float threshold(threshold) ;
		threshold:units = "K" ;
		threshold:standard_name = "air_temperature" ;
		threshold:spp__relative_to_threshold = "greater_than_or_equal_to" ;
	float projection_y_coordinate(projection_y_coordinate) ;
		projection_y_coordinate:axis = "Y" ;
		projection_y_coordinate:bounds = "projection_y_coordinate_bnds" ;
		projection_y_coordinate:units = "m" ;
		projection_y_coordinate:standard_name = "projection_y_coordinate" ;
	float projection_y_coordinate_bnds(projection_y_coordinate, bnds) ;
	float projection_x_coordinate(projection_x_coordinate) ;
		projection_x_coordinate:axis = "X" ;
		projection_x_coordinate:bounds = "projection_x_coordinate_bnds" ;
		projection_x_coordinate:units = "m" ;
		projection_x_coordinate:standard_name = "projection_x_coordinate" ;
	float projection_x_coordinate_bnds(projection_x_coordinate, bnds) ;
	int64 blend_time ;
		blend_time:units = "seconds since 1970-01-01 00:00:00" ;
		blend_time:long_name = "blend_time" ;
		blend_time:calendar = "gregorian" ;
	int forecast_period ;
		forecast_period:units = "seconds" ;
		forecast_period:standard_name = "forecast_period" ;
		forecast_period:deprecation_message = "forecast_period will be removed in future and should not be used" ;
	int64 forecast_reference_time ;
		forecast_reference_time:units = "seconds since 1970-01-01 00:00:00" ;
		forecast_reference_time:standard_name = "forecast_reference_time" ;
		forecast_reference_time:calendar = "gregorian" ;
		forecast_reference_time:deprecation_message = "forecast_reference_time will be removed in future and should not be used" ;
	float height ;
		height:units = "m" ;
		height:standard_name = "height" ;
		height:positive = "up" ;
	int64 time ;
		time:units = "seconds since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "gregorian" ;

// global attributes:
		:institution = "Met Office" ;
		:mosg__model_configuration = "gl_ens uk_ens" ;
		:source = "IMPROVER" ;
		:title = "IMPROVER Post-Processed Multi-Model Blend on UK 2 km Standard Grid" ;
		:Conventions = "CF-1.5" ;
data:

 threshold = 248.15, 253.15, 254.15, 255.15, 256.15, 257.15, 258.15, 259.15, 
    260.15, 261.15, 262.15, 263.15, 264.15, 265.15, 266.15, 267.15, 268.15, 
    269.15, 270.15, 271.15, 272.15, 273.15, 274.15, 275.15, 276.15, 277.15, 
    278.15, 279.15, 280.15, 281.15, 282.15, 283.15, 284.15, 285.15, 286.15, 
    287.15, 288.15, 289.15, 290.15, 291.15, 292.15, 293.15, 294.15, 295.15, 
    296.15, 297.15, 298.15, 299.15, 300.15, 301.15, 302.15, 303.15, 304.15, 
    305.15, 306.15, 307.15, 308.15, 309.15, 310.15, 311.15, 312.15, 313.15, 
    318.15 ;

 time = 1614960000 ;
}
