netcdf \20210315T0700Z-PT0001H00M-feels_like_temperature {
dimensions:
	percentile = 15 ;
	latitude = 960 ;
	longitude = 1280 ;
	bnds = 2 ;
variables:
	float feels_like_temperature(percentile, latitude, longitude) ;
		feels_like_temperature:long_name = "feels_like_temperature" ;
		feels_like_temperature:units = "K" ;
		feels_like_temperature:grid_mapping = "latitude_longitude" ;
		feels_like_temperature:coordinates = "blend_time forecast_period forecast_reference_time height time" ;
	int latitude_longitude ;
		latitude_longitude:grid_mapping_name = "latitude_longitude" ;
		latitude_longitude:longitude_of_prime_meridian = 0. ;
		latitude_longitude:earth_radius = 6371229. ;
	float percentile(percentile) ;
		percentile:units = "%" ;
		percentile:long_name = "percentile" ;
	float latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:bounds = "latitude_bnds" ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
	float latitude_bnds(latitude, bnds) ;
	float longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:bounds = "longitude_bnds" ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;
	float longitude_bnds(longitude, bnds) ;
	int64 blend_time ;
		blend_time:units = "seconds since 1970-01-01 00:00:00" ;
		blend_time:long_name = "blend_time" ;
		blend_time:calendar = "gregorian" ;
	int forecast_period ;
		forecast_period:units = "seconds" ;
		forecast_period:standard_name = "forecast_period" ;
		forecast_period:deprecation_message = "forecast_period will be removed in future and should not be used" ;
	int64 forecast_reference_time ;
		forecast_reference_time:units = "seconds since 1970-01-01 00:00:00" ;
		forecast_reference_time:standard_name = "forecast_reference_time" ;
		forecast_reference_time:calendar = "gregorian" ;
		forecast_reference_time:deprecation_message = "forecast_reference_time will be removed in future and should not be used" ;
	float height ;
		height:units = "m" ;
		height:standard_name = "height" ;
		height:positive = "up" ;
	int64 time ;
		time:units = "seconds since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "gregorian" ;

// global attributes:
		:institution = "Met Office" ;
		:mosg__model_configuration = "gl_ens" ;
		:source = "Met Office Unified Model" ;
		:title = "Post-Processed MOGREPS-G Model Forecast on Global 20 km Standard Grid" ;
		:Conventions = "CF-1.5" ;
data:

 percentile = 0, 5, 10, 20, 25, 30, 40, 50, 60, 70, 75, 80, 90, 95, 100 ;

 time = 1615791600 ;
}
