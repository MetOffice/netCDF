netcdf Fields_grid_conc_C1_T1_202505260100 {
dimensions:
	latitude = 261 ;
	longitude = 311 ;
	nbounds = 2 ;
	string23 = 23 ;
variables:
	float latitude(latitude) ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:axis = "Y" ;
		latitude:valid_min = 48.f ;
		latitude:valid_max = 61.f ;
		latitude:bounds = "latitude_bounds" ;
	float longitude(longitude) ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:axis = "X" ;
		longitude:valid_min = -11.f ;
		longitude:valid_max = 4.5f ;
		longitude:bounds = "longitude_bounds" ;
	float latitude_bounds(latitude, nbounds) ;
		latitude_bounds:comment = "Bounds" ;
	float longitude_bounds(longitude, nbounds) ;
		longitude_bounds:comment = "Bounds" ;
	int time_0 ;
		time_0:standard_name = "time" ;
		time_0:long_name = "time" ;
		time_0:units = "minutes since 1970-01-01 00:00:00" ;
		time_0:calendar = "gregorian" ;
		time_0:bounds = "time_bnds_0" ;
	int time_bnds_0(nbounds) ;
		time_bnds_0:long_name = "start_and_end_point" ;
	int forecast_reference_time ;
		forecast_reference_time:standard_name = "forecast_reference_time" ;
		forecast_reference_time:long_name = "forecast_reference_time" ;
		forecast_reference_time:units = "minutes since 1970-01-01 00:00:00" ;
		forecast_reference_time:calendar = "gregorian" ;
	int latitude_longitude ;
		latitude_longitude:grid_mapping_name = "latitude_longitude" ;
		latitude_longitude:longitude_of_prime_meridian = 0.f ;
		latitude_longitude:earth_radius = 6371229.f ;
	float height ;
		height:standard_name = "height" ;
		height:comment = "height above ground level" ;
		height:units = "m" ;
		height:long_name = "height above ground level" ;
		height:axis = "Z" ;
		height:positive = "up" ;
		height:reference_datum = "ground level" ;
		height:bounds = "height_bnds" ;
	float height_bnds(nbounds) ;
		height_bnds:long_name = "height above ground level start and end point" ;
	float GRASS_POLLEN_CONCENTRATION(latitude, longitude) ;
		GRASS_POLLEN_CONCENTRATION:long_name = "GRASS_POLLEN_CONCENTRATION" ;
		GRASS_POLLEN_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		GRASS_POLLEN_CONCENTRATION:field_name = "Unnamed Field Req 2" ;
		GRASS_POLLEN_CONCENTRATION:units = "g / m^3" ;
		GRASS_POLLEN_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		GRASS_POLLEN_CONCENTRATION:quantity = "Concentration" ;
		GRASS_POLLEN_CONCENTRATION:species = "GRASS_POLLEN" ;
		GRASS_POLLEN_CONCENTRATION:species_category = "POLLEN" ;
		GRASS_POLLEN_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		GRASS_POLLEN_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		GRASS_POLLEN_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		GRASS_POLLEN_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float BIRCH_POLLEN_CONCENTRATION(latitude, longitude) ;
		BIRCH_POLLEN_CONCENTRATION:long_name = "BIRCH_POLLEN_CONCENTRATION" ;
		BIRCH_POLLEN_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		BIRCH_POLLEN_CONCENTRATION:field_name = "Unnamed Field Req 6" ;
		BIRCH_POLLEN_CONCENTRATION:units = "g / m^3" ;
		BIRCH_POLLEN_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		BIRCH_POLLEN_CONCENTRATION:quantity = "Concentration" ;
		BIRCH_POLLEN_CONCENTRATION:species = "BIRCH_POLLEN" ;
		BIRCH_POLLEN_CONCENTRATION:species_category = "POLLEN" ;
		BIRCH_POLLEN_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		BIRCH_POLLEN_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		BIRCH_POLLEN_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		BIRCH_POLLEN_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float OAK_POLLEN_CONCENTRATION(latitude, longitude) ;
		OAK_POLLEN_CONCENTRATION:long_name = "OAK_POLLEN_CONCENTRATION" ;
		OAK_POLLEN_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		OAK_POLLEN_CONCENTRATION:field_name = "Unnamed Field Req 10" ;
		OAK_POLLEN_CONCENTRATION:units = "g / m^3" ;
		OAK_POLLEN_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		OAK_POLLEN_CONCENTRATION:quantity = "Concentration" ;
		OAK_POLLEN_CONCENTRATION:species = "OAK_POLLEN" ;
		OAK_POLLEN_CONCENTRATION:species_category = "POLLEN" ;
		OAK_POLLEN_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		OAK_POLLEN_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		OAK_POLLEN_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		OAK_POLLEN_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float ALDER_POLLEN_CONCENTRATION(latitude, longitude) ;
		ALDER_POLLEN_CONCENTRATION:long_name = "ALDER_POLLEN_CONCENTRATION" ;
		ALDER_POLLEN_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		ALDER_POLLEN_CONCENTRATION:field_name = "Unnamed Field Req 14" ;
		ALDER_POLLEN_CONCENTRATION:units = "g / m^3" ;
		ALDER_POLLEN_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		ALDER_POLLEN_CONCENTRATION:quantity = "Concentration" ;
		ALDER_POLLEN_CONCENTRATION:species = "ALDER_POLLEN" ;
		ALDER_POLLEN_CONCENTRATION:species_category = "POLLEN" ;
		ALDER_POLLEN_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		ALDER_POLLEN_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		ALDER_POLLEN_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		ALDER_POLLEN_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float HAZEL_POLLEN_CONCENTRATION(latitude, longitude) ;
		HAZEL_POLLEN_CONCENTRATION:long_name = "HAZEL_POLLEN_CONCENTRATION" ;
		HAZEL_POLLEN_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		HAZEL_POLLEN_CONCENTRATION:field_name = "Unnamed Field Req 18" ;
		HAZEL_POLLEN_CONCENTRATION:units = "g / m^3" ;
		HAZEL_POLLEN_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		HAZEL_POLLEN_CONCENTRATION:quantity = "Concentration" ;
		HAZEL_POLLEN_CONCENTRATION:species = "HAZEL_POLLEN" ;
		HAZEL_POLLEN_CONCENTRATION:species_category = "POLLEN" ;
		HAZEL_POLLEN_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		HAZEL_POLLEN_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		HAZEL_POLLEN_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		HAZEL_POLLEN_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float NETTLE_POLLEN_CONCENTRATION(latitude, longitude) ;
		NETTLE_POLLEN_CONCENTRATION:long_name = "NETTLE_POLLEN_CONCENTRATION" ;
		NETTLE_POLLEN_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		NETTLE_POLLEN_CONCENTRATION:field_name = "Unnamed Field Req 22" ;
		NETTLE_POLLEN_CONCENTRATION:units = "g / m^3" ;
		NETTLE_POLLEN_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		NETTLE_POLLEN_CONCENTRATION:quantity = "Concentration" ;
		NETTLE_POLLEN_CONCENTRATION:species = "NETTLE_POLLEN" ;
		NETTLE_POLLEN_CONCENTRATION:species_category = "POLLEN" ;
		NETTLE_POLLEN_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		NETTLE_POLLEN_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		NETTLE_POLLEN_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		NETTLE_POLLEN_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float ASH_POLLEN_CONCENTRATION(latitude, longitude) ;
		ASH_POLLEN_CONCENTRATION:long_name = "ASH_POLLEN_CONCENTRATION" ;
		ASH_POLLEN_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		ASH_POLLEN_CONCENTRATION:field_name = "Unnamed Field Req 26" ;
		ASH_POLLEN_CONCENTRATION:units = "g / m^3" ;
		ASH_POLLEN_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		ASH_POLLEN_CONCENTRATION:quantity = "Concentration" ;
		ASH_POLLEN_CONCENTRATION:species = "ASH_POLLEN" ;
		ASH_POLLEN_CONCENTRATION:species_category = "POLLEN" ;
		ASH_POLLEN_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		ASH_POLLEN_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		ASH_POLLEN_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		ASH_POLLEN_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float PLANE_POLLEN_CONCENTRATION(latitude, longitude) ;
		PLANE_POLLEN_CONCENTRATION:long_name = "PLANE_POLLEN_CONCENTRATION" ;
		PLANE_POLLEN_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		PLANE_POLLEN_CONCENTRATION:field_name = "Unnamed Field Req 30" ;
		PLANE_POLLEN_CONCENTRATION:units = "g / m^3" ;
		PLANE_POLLEN_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		PLANE_POLLEN_CONCENTRATION:quantity = "Concentration" ;
		PLANE_POLLEN_CONCENTRATION:species = "PLANE_POLLEN" ;
		PLANE_POLLEN_CONCENTRATION:species_category = "POLLEN" ;
		PLANE_POLLEN_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		PLANE_POLLEN_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		PLANE_POLLEN_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		PLANE_POLLEN_CONCENTRATION:cell_methods = "time: mean height: mean" ;

// global attributes:
		:title = "Pollen_test" ;
		:Conventions = "CF-1.8" ;
		:history = "NAME 13/11/2025 15:39:31.175 UTC" ;
		:source = "Met Office NAME model" ;
		:institution = "NA" ;
		:reference = "https://doi.org/10.1007/978-0-387-68854-1_62" ;
		:comment = "none" ;
		:name_version = "NAME III (development version 8.7+)" ;
		:run_time = "13/11/2025 15:39:31.175 UTC" ;
		:run_duration = "12hr 0min" ;
		:met_data = "NWP Flow.UKV_PT1_flow; NWP Flow.UKV_PT2_flow; NWP Flow.UKV_PT3_flow; NWP Flow.UKV_PT4_flow; NWP Flow.UKV_PT5_flow; NWP Flow.UKV_PT6_flow; NWP Flow.UKV_PT7_flow; NWP Flow.UKV_PT8_flow; NWP Flow.UKV_PT9_flow; NWP Flow.UKV_PT10_flow; NWP Flow.UKV_PT11_flow; NWP Flow.UKV_PT12_flow; NWP Flow.UKV_PT13_flow; NWP Flow.UKV_PT14_flow; NWP Flow.UKV_PT15_flow; NWP Flow.UKV_PT16_flow; NWP Flow.Regional" ;
		:name_netcdf_out_vers = "0.1" ;
		:start_of_release = "-infinity" ;
		:end_of_release = "infinity" ;
		:source_strength = "Multiple Sources" ;
		:release_location = "Multiple Sources" ;
		:release_height = "Multiple Sources" ;
}
