netcdf \20210326T0000Z-PT0000H00M-soil_temperature_on_soil_levels {
dimensions:
	depth = 4 ;
	latitude = 1920 ;
	longitude = 2560 ;
	bnds = 2 ;
variables:
	float soil_temperature(depth, latitude, longitude) ;
		soil_temperature:_FillValue = NaNf ;
		soil_temperature:least_significant_digit = 1LL ;
		soil_temperature:standard_name = "soil_temperature" ;
		soil_temperature:units = "K" ;
		soil_temperature:grid_mapping = "latitude_longitude" ;
		soil_temperature:coordinates = "forecast_period forecast_reference_time time" ;
	int latitude_longitude ;
		latitude_longitude:grid_mapping_name = "latitude_longitude" ;
		latitude_longitude:longitude_of_prime_meridian = 0. ;
		latitude_longitude:earth_radius = 6371229. ;
	float depth(depth) ;
		depth:axis = "Z" ;
		depth:bounds = "depth_bnds" ;
		depth:units = "m" ;
		depth:standard_name = "depth" ;
		depth:positive = "down" ;
	float depth_bnds(depth, bnds) ;
	float latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:bounds = "latitude_bnds" ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
	float latitude_bnds(latitude, bnds) ;
	float longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:bounds = "longitude_bnds" ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;
	float longitude_bnds(longitude, bnds) ;
	int forecast_period ;
		forecast_period:units = "seconds" ;
		forecast_period:standard_name = "forecast_period" ;
	int64 forecast_reference_time ;
		forecast_reference_time:units = "seconds since 1970-01-01 00:00:00" ;
		forecast_reference_time:standard_name = "forecast_reference_time" ;
		forecast_reference_time:calendar = "gregorian" ;
	int64 time ;
		time:units = "seconds since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "gregorian" ;

// global attributes:
		:history = "2021-03-26T04:09:12Z: StaGE Decoupler" ;
		:institution = "Met Office" ;
		:mosg__forecast_run_duration = "PT168H" ;
		:mosg__grid_domain = "global" ;
		:mosg__grid_type = "standard" ;
		:mosg__grid_version = "1.6.0" ;
		:mosg__model_configuration = "gl_det" ;
		:source = "Met Office Unified Model" ;
		:title = "Global Model Forecast on Global 10 km Standard Grid" ;
		:um_version = "11.5" ;
		:Conventions = "CF-1.7, UKMO-1.0" ;
data:

 time = 1616716800 ;
}
