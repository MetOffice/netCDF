netcdf Fields_grid2_C1_T1_201807031200 {
dimensions:
	latitude = 200 ;
	longitude = 200 ;
	nbounds = 2 ;
	string23 = 23 ;
variables:
	float latitude(latitude) ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:axis = "Y" ;
		latitude:valid_min = 51.39275f ;
		latitude:valid_max = 51.61164f ;
		latitude:bounds = "latitude_bounds" ;
	float longitude(longitude) ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:axis = "X" ;
		longitude:valid_min = -0.306088f ;
		longitude:valid_max = 0.05211202f ;
		longitude:bounds = "longitude_bounds" ;
	float latitude_bounds(latitude, nbounds) ;
		latitude_bounds:comment = "Bounds" ;
	float longitude_bounds(longitude, nbounds) ;
		longitude_bounds:comment = "Bounds" ;
	int time_0 ;
		time_0:standard_name = "time" ;
		time_0:long_name = "time" ;
		time_0:units = "minutes since 1970-01-01 00:00:00" ;
		time_0:calendar = "gregorian" ;
		time_0:bounds = "time_bnds_0" ;
	int time_bnds_0(nbounds) ;
		time_bnds_0:long_name = "start_and_end_point" ;
	int forecast_reference_time ;
		forecast_reference_time:standard_name = "forecast_reference_time" ;
		forecast_reference_time:long_name = "forecast_reference_time" ;
		forecast_reference_time:units = "minutes since 1970-01-01 00:00:00" ;
		forecast_reference_time:calendar = "gregorian" ;
	int latitude_longitude ;
		latitude_longitude:grid_mapping_name = "latitude_longitude" ;
		latitude_longitude:longitude_of_prime_meridian = 0.f ;
		latitude_longitude:earth_radius = 6371229.f ;
	float height ;
		height:standard_name = "height" ;
		height:comment = "height above ground level" ;
		height:units = "m" ;
		height:long_name = "height above ground level" ;
		height:axis = "Z" ;
		height:positive = "up" ;
		height:reference_datum = "ground level" ;
		height:bounds = "height_bnds" ;
	float height_bnds(nbounds) ;
		height_bnds:long_name = "height above ground level start and end point" ;
	float TRACER_AIR_CONCENTRATION(latitude, longitude) ;
		TRACER_AIR_CONCENTRATION:long_name = "TRACER_AIR_CONCENTRATION" ;
		TRACER_AIR_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		TRACER_AIR_CONCENTRATION:field_name = "Unnamed Field Req 1" ;
		TRACER_AIR_CONCENTRATION:units = "g / m^3" ;
		TRACER_AIR_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		TRACER_AIR_CONCENTRATION:quantity = "Air Concentration" ;
		TRACER_AIR_CONCENTRATION:source_or_sourcegroup = "All sources" ;
		TRACER_AIR_CONCENTRATION:species = "TRACER" ;
		TRACER_AIR_CONCENTRATION:species_category = "CHEMISTRY-SPECIES" ;
		TRACER_AIR_CONCENTRATION:time_av_int_info = "3hr 0min average" ;
		TRACER_AIR_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		TRACER_AIR_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		TRACER_AIR_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float TRACER_WET_DEPOSITION(latitude, longitude) ;
		TRACER_WET_DEPOSITION:long_name = "TRACER_WET_DEPOSITION" ;
		TRACER_WET_DEPOSITION:grid_mapping = "latitude_longitude" ;
		TRACER_WET_DEPOSITION:field_name = "Unnamed Field Req 3" ;
		TRACER_WET_DEPOSITION:units = "g / m^2" ;
		TRACER_WET_DEPOSITION:coordinates = "time_0 forecast_reference_time" ;
		TRACER_WET_DEPOSITION:quantity = "Wet Deposition" ;
		TRACER_WET_DEPOSITION:source_or_sourcegroup = "All sources" ;
		TRACER_WET_DEPOSITION:species = "TRACER" ;
		TRACER_WET_DEPOSITION:species_category = "CHEMISTRY-SPECIES" ;
		TRACER_WET_DEPOSITION:time_av_int_info = "3hr 0min integral" ;
		TRACER_WET_DEPOSITION:horizontal_av_int_info = "No horizontal averaging" ;
		TRACER_WET_DEPOSITION:cell_methods = "time: sum" ;
	float TRACER_DRY_DEPOSITION(latitude, longitude) ;
		TRACER_DRY_DEPOSITION:long_name = "TRACER_DRY_DEPOSITION" ;
		TRACER_DRY_DEPOSITION:grid_mapping = "latitude_longitude" ;
		TRACER_DRY_DEPOSITION:field_name = "Unnamed Field Req 4" ;
		TRACER_DRY_DEPOSITION:units = "g / m^2" ;
		TRACER_DRY_DEPOSITION:coordinates = "time_0 forecast_reference_time" ;
		TRACER_DRY_DEPOSITION:quantity = "Dry Deposition" ;
		TRACER_DRY_DEPOSITION:source_or_sourcegroup = "All sources" ;
		TRACER_DRY_DEPOSITION:species = "TRACER" ;
		TRACER_DRY_DEPOSITION:species_category = "CHEMISTRY-SPECIES" ;
		TRACER_DRY_DEPOSITION:time_av_int_info = "3hr 0min integral" ;
		TRACER_DRY_DEPOSITION:horizontal_av_int_info = "No horizontal averaging" ;
		TRACER_DRY_DEPOSITION:cell_methods = "time: sum" ;
	float TRACER_DEPOSITION(latitude, longitude) ;
		TRACER_DEPOSITION:long_name = "TRACER_DEPOSITION" ;
		TRACER_DEPOSITION:grid_mapping = "latitude_longitude" ;
		TRACER_DEPOSITION:field_name = "Unnamed Field Req 5" ;
		TRACER_DEPOSITION:units = "g / m^2" ;
		TRACER_DEPOSITION:coordinates = "time_0 forecast_reference_time" ;
		TRACER_DEPOSITION:quantity = "Deposition" ;
		TRACER_DEPOSITION:source_or_sourcegroup = "All sources" ;
		TRACER_DEPOSITION:species = "TRACER" ;
		TRACER_DEPOSITION:species_category = "CHEMISTRY-SPECIES" ;
		TRACER_DEPOSITION:time_av_int_info = "3hr 0min integral" ;
		TRACER_DEPOSITION:horizontal_av_int_info = "No horizontal averaging" ;
		TRACER_DEPOSITION:cell_methods = "time: sum" ;

// global attributes:
		:title = "Operational - CHEMET Test 1" ;
		:Conventions = "CF-1.8" ;
		:history = "NAME 13/11/2025 15:39:18.386 UTC" ;
		:source = "Met Office NAME model" ;
		:institution = "NA" ;
		:reference = "https://doi.org/10.1007/978-0-387-68854-1_62" ;
		:comment = "none" ;
		:name_version = "NAME III (development version 8.7+)" ;
		:run_time = "13/11/2025 15:39:18.386 UTC" ;
		:run_duration = "3hr 0min" ;
		:met_data = "NWP Flow.UKV_PT1_flow; NWP Flow.UKV_PT2_flow; NWP Flow.UKV_PT3_flow; NWP Flow.UKV_PT4_flow; NWP Flow.UKV_PT5_flow; NWP Flow.UKV_PT6_flow; NWP Flow.UKV_PT7_flow; NWP Flow.UKV_PT8_flow; NWP Flow.UKV_PT9_flow; NWP Flow.UKV_PT10_flow; NWP Flow.UKV_PT11_flow; NWP Flow.UKV_PT12_flow; NWP Flow.UKV_PT13_flow; NWP Flow.UKV_PT14_flow; NWP Flow.UKV_PT15_flow; NWP Flow.UKV_PT16_flow; NWP Flow.Global_PT2_flow" ;
		:name_netcdf_out_vers = "0.1" ;
		:start_of_release = "03/07/2018 09:00 UTC" ;
		:end_of_release = "03/07/2018 12:00 UTC" ;
		:source_strength = "1 g/s" ;
		:release_location = "0.1270W   51.5022N" ;
		:release_height = "0.000 to 10.000m agl" ;
}
