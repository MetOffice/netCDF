netcdf QVA_grid1_C1_T1_201810221200 {
dimensions:
	latitude = 720 ;
	longitude = 1440 ;
	nbounds = 2 ;
	string23 = 23 ;
	flight_level = 12 ;
variables:
	float latitude(latitude) ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:axis = "Y" ;
		latitude:valid_min = -89.875f ;
		latitude:valid_max = 89.875f ;
		latitude:bounds = "latitude_bounds" ;
	float longitude(longitude) ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:axis = "X" ;
		longitude:valid_min = -179.875f ;
		longitude:valid_max = 179.875f ;
		longitude:bounds = "longitude_bounds" ;
	float latitude_bounds(latitude, nbounds) ;
		latitude_bounds:comment = "Bounds" ;
	float longitude_bounds(longitude, nbounds) ;
		longitude_bounds:comment = "Bounds" ;
	float flight_level(flight_level) ;
		flight_level:units = "geopotential hft" ;
		flight_level:long_name = "flight level" ;
		flight_level:axis = "Z" ;
		flight_level:positive = "up" ;
		flight_level:valid_min = 25.f ;
		flight_level:valid_max = 575.f ;
		flight_level:bounds = "flight_level_bounds" ;
		flight_level:reference_datum = "sea level pressure datum of 1013.25 hPa" ;
	float flight_level_bounds(flight_level, nbounds) ;
		flight_level_bounds:comment = "for each level, lower and upper bounds" ;
	int time_0 ;
		time_0:standard_name = "time" ;
		time_0:long_name = "time" ;
		time_0:units = "minutes since 1970-01-01 00:00:00" ;
		time_0:calendar = "gregorian" ;
		time_0:bounds = "time_bnds_0" ;
	int time_bnds_0(nbounds) ;
		time_bnds_0:long_name = "start_and_end_point" ;
	int forecast_reference_time ;
		forecast_reference_time:standard_name = "forecast_reference_time" ;
		forecast_reference_time:long_name = "forecast_reference_time" ;
		forecast_reference_time:units = "minutes since 1970-01-01 00:00:00" ;
		forecast_reference_time:calendar = "gregorian" ;
	int latitude_longitude ;
		latitude_longitude:grid_mapping_name = "latitude_longitude" ;
		latitude_longitude:longitude_of_prime_meridian = 0.f ;
		latitude_longitude:earth_radius = 6371229.f ;
	float VOLCANIC_ASH_AIR_CONCENTRATION(flight_level, latitude, longitude) ;
		VOLCANIC_ASH_AIR_CONCENTRATION:long_name = "VOLCANIC_ASH_AIR_CONCENTRATION" ;
		VOLCANIC_ASH_AIR_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		VOLCANIC_ASH_AIR_CONCENTRATION:field_name = "Unnamed Field Req 1" ;
		VOLCANIC_ASH_AIR_CONCENTRATION:units = "g / m^3" ;
		VOLCANIC_ASH_AIR_CONCENTRATION:coordinates = "time_0 forecast_reference_time" ;
		VOLCANIC_ASH_AIR_CONCENTRATION:quantity = "Air Concentration" ;
		VOLCANIC_ASH_AIR_CONCENTRATION:source_or_sourcegroup = "All sources" ;
		VOLCANIC_ASH_AIR_CONCENTRATION:species = "VOLCANIC_ASH" ;
		VOLCANIC_ASH_AIR_CONCENTRATION:species_category = "VOLCANIC" ;
		VOLCANIC_ASH_AIR_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		VOLCANIC_ASH_AIR_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		VOLCANIC_ASH_AIR_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		VOLCANIC_ASH_AIR_CONCENTRATION:cell_methods = "time: mean flight_level: mean" ;

// global attributes:
		:title = "Operational - VAAC UM Global" ;
		:Conventions = "CF-1.8" ;
		:history = "NAME 13/11/2025 15:44:58.959 UTC" ;
		:source = "Met Office NAME model" ;
		:institution = "NA" ;
		:reference = "https://doi.org/10.1007/978-0-387-68854-1_62" ;
		:comment = "none" ;
		:name_version = "NAME III (development version 8.7+)" ;
		:run_time = "13/11/2025 15:44:58.959 UTC" ;
		:run_duration = "11day 12hr 10min" ;
		:met_data = "NWP Flow.Global_PT1_flow; NWP Flow.Global_PT2_flow; NWP Flow.Global_PT3_flow; NWP Flow.Global_PT4_flow; NWP Flow.Global_PT5_flow; NWP Flow.Global_PT6_flow; NWP Flow.Global_PT7_flow; NWP Flow.Global_PT8_flow; NWP Flow.Global_PT9_flow; NWP Flow.Global_PT10_flow; NWP Flow.Global_PT11_flow; NWP Flow.Global_PT12_flow; NWP Flow.Global_PT13_flow; NWP Flow.Global_PT14_flow" ;
		:name_netcdf_out_vers = "0.1" ;
		:start_of_release = "22/10/2018 09:45 UTC" ;
		:end_of_release = "30/06/2028 00:00 UTC" ;
		:source_strength = "4.697695E+07 g/s" ;
		:release_location = "19.6300W   63.6300N" ;
		:release_height = "5825.500m asl +/- 4174.500m" ;
}
