netcdf Fields_grid1_C1_T1_201807040000 {
dimensions:
	latitude = 480 ;
	longitude = 640 ;
	nbounds = 2 ;
	string23 = 23 ;
variables:
	float latitude(latitude) ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:axis = "Y" ;
		latitude:valid_min = -89.8125f ;
		latitude:valid_max = 89.8125f ;
		latitude:bounds = "latitude_bounds" ;
	float longitude(longitude) ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:axis = "X" ;
		longitude:valid_min = 0.28125f ;
		longitude:valid_max = 359.7188f ;
		longitude:bounds = "longitude_bounds" ;
	float latitude_bounds(latitude, nbounds) ;
		latitude_bounds:comment = "Bounds" ;
	float longitude_bounds(longitude, nbounds) ;
		longitude_bounds:comment = "Bounds" ;
	int time_0 ;
		time_0:standard_name = "time" ;
		time_0:long_name = "time" ;
		time_0:units = "minutes since 1970-01-01 00:00:00" ;
		time_0:calendar = "gregorian" ;
		time_0:bounds = "time_bnds_0" ;
	int time_bnds_0(nbounds) ;
		time_bnds_0:long_name = "start_and_end_point" ;
	int time_1 ;
		time_1:standard_name = "time" ;
		time_1:long_name = "time" ;
		time_1:units = "minutes since 1970-01-01 00:00:00" ;
		time_1:calendar = "gregorian" ;
		time_1:bounds = "time_bnds_1" ;
	int time_bnds_1(nbounds) ;
		time_bnds_1:long_name = "start_and_end_point" ;
	int forecast_reference_time ;
		forecast_reference_time:standard_name = "forecast_reference_time" ;
		forecast_reference_time:long_name = "forecast_reference_time" ;
		forecast_reference_time:units = "minutes since 1970-01-01 00:00:00" ;
		forecast_reference_time:calendar = "gregorian" ;
	int latitude_longitude ;
		latitude_longitude:grid_mapping_name = "latitude_longitude" ;
		latitude_longitude:longitude_of_prime_meridian = 0.f ;
		latitude_longitude:earth_radius = 6371229.f ;
	float height ;
		height:standard_name = "height" ;
		height:comment = "height above ground level" ;
		height:units = "m" ;
		height:long_name = "height above ground level" ;
		height:axis = "Z" ;
		height:positive = "up" ;
		height:reference_datum = "ground level" ;
		height:bounds = "height_bnds" ;
	float height_bnds(nbounds) ;
		height_bnds:long_name = "height above ground level start and end point" ;
	float CAESIUM_137_AIR_CONCENTRATION(latitude, longitude) ;
		CAESIUM_137_AIR_CONCENTRATION:long_name = "CAESIUM_137_AIR_CONCENTRATION" ;
		CAESIUM_137_AIR_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		CAESIUM_137_AIR_CONCENTRATION:field_name = "Unnamed Field Req 1" ;
		CAESIUM_137_AIR_CONCENTRATION:units = "Bq s / m^3" ;
		CAESIUM_137_AIR_CONCENTRATION:coordinates = "time_1 forecast_reference_time height" ;
		CAESIUM_137_AIR_CONCENTRATION:quantity = "Air Concentration" ;
		CAESIUM_137_AIR_CONCENTRATION:source_or_sourcegroup = "All sources" ;
		CAESIUM_137_AIR_CONCENTRATION:species = "CAESIUM-137" ;
		CAESIUM_137_AIR_CONCENTRATION:species_category = "RADIONUCLIDE" ;
		CAESIUM_137_AIR_CONCENTRATION:time_av_int_info = "1day 0hr 0min integral" ;
		CAESIUM_137_AIR_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		CAESIUM_137_AIR_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		CAESIUM_137_AIR_CONCENTRATION:cell_methods = "time: sum height: mean" ;
	float CAESIUM_137_DEPOSITION(latitude, longitude) ;
		CAESIUM_137_DEPOSITION:long_name = "CAESIUM_137_DEPOSITION" ;
		CAESIUM_137_DEPOSITION:grid_mapping = "latitude_longitude" ;
		CAESIUM_137_DEPOSITION:field_name = "Unnamed Field Req 2" ;
		CAESIUM_137_DEPOSITION:units = "Bq / m^2" ;
		CAESIUM_137_DEPOSITION:coordinates = "time_0 forecast_reference_time" ;
		CAESIUM_137_DEPOSITION:quantity = "Deposition" ;
		CAESIUM_137_DEPOSITION:source_or_sourcegroup = "All sources" ;
		CAESIUM_137_DEPOSITION:species = "CAESIUM-137" ;
		CAESIUM_137_DEPOSITION:species_category = "RADIONUCLIDE" ;
		CAESIUM_137_DEPOSITION:time_av_int_info = "3day 0hr 0min integral" ;
		CAESIUM_137_DEPOSITION:horizontal_av_int_info = "No horizontal averaging" ;
		CAESIUM_137_DEPOSITION:cell_methods = "time: sum" ;

// global attributes:
		:title = "Operational - RSMC Test 1" ;
		:Conventions = "CF-1.8" ;
		:history = "NAME 13/11/2025 15:39:35.444 UTC" ;
		:source = "Met Office NAME model" ;
		:institution = "NA" ;
		:reference = "https://doi.org/10.1007/978-0-387-68854-1_62" ;
		:comment = "none" ;
		:name_version = "NAME III (development version 8.7+)" ;
		:run_time = "13/11/2025 15:39:35.444 UTC" ;
		:run_duration = "3day 0hr 0min" ;
		:met_data = "NWP Flow.Global_PT1_flow; NWP Flow.Global_PT2_flow; NWP Flow.Global_PT3_flow; NWP Flow.Global_PT4_flow; NWP Flow.Global_PT5_flow; NWP Flow.Global_PT6_flow; NWP Flow.Global_PT7_flow; NWP Flow.Global_PT8_flow; NWP Flow.Global_PT9_flow; NWP Flow.Global_PT10_flow; NWP Flow.Global_PT11_flow; NWP Flow.Global_PT12_flow; NWP Flow.Global_PT13_flow; NWP Flow.Global_PT14_flow" ;
		:name_netcdf_out_vers = "0.1" ;
		:start_of_release = "03/07/2018 10:00 UTC" ;
		:end_of_release = "03/07/2018 16:00 UTC" ;
		:source_strength = "4.630556E-05 Bq/s" ;
		:release_location = "30.0991E   51.3896N" ;
		:release_height = "0.000 to 500.000m agl" ;
}
