netcdf NonSpatialDimensions {
dimensions:
	axis_nbounds = 2 ;
	Two = 2 ;
	nMesh2d_face_node = 56 ;
	nMesh2d_face_edge = 108 ;
	nMesh2d_face_face = 54 ;
	nMesh2d_face_vertex = 4 ;
	mutable_categories = 3 ;
	str_len = 255 ;
	mutable_numbers = 2 ;
	immutable_categories = 3 ;
	immutable_numbers = 3 ;
	time_counter = UNLIMITED ; // (5 currently)
variables:
	int Mesh2d_face ;
		Mesh2d_face:cf_role = "mesh_topology" ;
		Mesh2d_face:long_name = "Topology data of 2D unstructured mesh" ;
		Mesh2d_face:topology_dimension = 2 ;
		Mesh2d_face:node_coordinates = "Mesh2d_face_node_x Mesh2d_face_node_y" ;
		Mesh2d_face:edge_coordinates = "Mesh2d_face_edge_x Mesh2d_face_edge_y" ;
		Mesh2d_face:edge_node_connectivity = "Mesh2d_face_edge_nodes" ;
		Mesh2d_face:face_coordinates = "Mesh2d_face_face_x Mesh2d_face_face_y" ;
		Mesh2d_face:face_node_connectivity = "Mesh2d_face_face_nodes" ;
	float Mesh2d_face_node_x(nMesh2d_face_node) ;
		Mesh2d_face_node_x:standard_name = "longitude" ;
		Mesh2d_face_node_x:long_name = "Longitude of mesh nodes." ;
		Mesh2d_face_node_x:units = "degrees_east" ;
	float Mesh2d_face_node_y(nMesh2d_face_node) ;
		Mesh2d_face_node_y:standard_name = "latitude" ;
		Mesh2d_face_node_y:long_name = "Latitude of mesh nodes." ;
		Mesh2d_face_node_y:units = "degrees_north" ;
	float Mesh2d_face_edge_x(nMesh2d_face_edge) ;
		Mesh2d_face_edge_x:standard_name = "longitude" ;
		Mesh2d_face_edge_x:long_name = "Characteristic longitude of mesh edges." ;
		Mesh2d_face_edge_x:units = "degrees_east" ;
	float Mesh2d_face_edge_y(nMesh2d_face_edge) ;
		Mesh2d_face_edge_y:standard_name = "latitude" ;
		Mesh2d_face_edge_y:long_name = "Characteristic latitude of mesh edges." ;
		Mesh2d_face_edge_y:units = "degrees_north" ;
	int Mesh2d_face_edge_nodes(nMesh2d_face_edge, Two) ;
		Mesh2d_face_edge_nodes:cf_role = "edge_node_connectivity" ;
		Mesh2d_face_edge_nodes:long_name = "Maps every edge/link to two nodes that it connects." ;
		Mesh2d_face_edge_nodes:start_index = 0 ;
	float Mesh2d_face_face_x(nMesh2d_face_face) ;
		Mesh2d_face_face_x:standard_name = "longitude" ;
		Mesh2d_face_face_x:long_name = "Characteristic longitude of mesh faces." ;
		Mesh2d_face_face_x:units = "degrees_east" ;
	float Mesh2d_face_face_y(nMesh2d_face_face) ;
		Mesh2d_face_face_y:standard_name = "latitude" ;
		Mesh2d_face_face_y:long_name = "Characteristic latitude of mesh faces." ;
		Mesh2d_face_face_y:units = "degrees_north" ;
	int Mesh2d_face_face_nodes(nMesh2d_face_face, nMesh2d_face_vertex) ;
		Mesh2d_face_face_nodes:cf_role = "face_node_connectivity" ;
		Mesh2d_face_face_nodes:long_name = "Maps every face to its corner nodes." ;
		Mesh2d_face_face_nodes:start_index = 0 ;
	int Mesh2d_face_face_edges(nMesh2d_face_face, nMesh2d_face_vertex) ;
		Mesh2d_face_face_edges:cf_role = "face_edge_connectivity" ;
		Mesh2d_face_face_edges:long_name = "Maps every face to its edges." ;
		Mesh2d_face_face_edges:start_index = 0 ;
		Mesh2d_face_face_edges:_FillValue = 999999 ;
	int Mesh2d_face_edge_face_links(nMesh2d_face_edge, Two) ;
		Mesh2d_face_edge_face_links:cf_role = "edge_face connectivity" ;
		Mesh2d_face_edge_face_links:long_name = "neighbor faces for edges" ;
		Mesh2d_face_edge_face_links:start_index = 0 ;
		Mesh2d_face_edge_face_links:_FillValue = -999 ;
		Mesh2d_face_edge_face_links:comment = "missing neighbor faces are indicated using _FillValue" ;
	int Mesh2d_face_face_links(nMesh2d_face_face, nMesh2d_face_vertex) ;
		Mesh2d_face_face_links:cf_role = "face_face connectivity" ;
		Mesh2d_face_face_links:long_name = "Indicates which other faces neighbor each face" ;
		Mesh2d_face_face_links:start_index = 0 ;
		Mesh2d_face_face_links:_FillValue = 999999 ;
		Mesh2d_face_face_links:flag_values = -1 ;
		Mesh2d_face_face_links:flag_meanings = "out_of_mesh" ;
	char mutable_categories(mutable_categories, str_len) ;
		mutable_categories:name = "mutable_categories" ;
	char mutable_numbers(mutable_numbers, str_len) ;
		mutable_numbers:name = "mutable_numbers" ;
		mutable_numbers:units = "other units" ;
	char immutable_categories(immutable_categories, str_len) ;
		immutable_categories:name = "immutable_categories" ;
	char immutable_numbers(immutable_numbers, str_len) ;
		immutable_numbers:name = "immutable_numbers" ;
		immutable_numbers:units = "other units" ;
	double time_instant(time_counter) ;
		time_instant:standard_name = "time" ;
		time_instant:long_name = "Time axis" ;
		time_instant:calendar = "gregorian" ;
		time_instant:units = "seconds since 0000-01-01 00:00:00" ;
		time_instant:time_origin = "0000-01-01 00:00:00" ;
		time_instant:bounds = "time_instant_bounds" ;
	double time_instant_bounds(time_counter, axis_nbounds) ;
	double colours__mutable_categories__instant_1ts(time_counter, mutable_categories, nMesh2d_face_face) ;
		colours__mutable_categories__instant_1ts:standard_name = "mutable_categories" ;
		colours__mutable_categories__instant_1ts:units = "arbitrary units" ;
		colours__mutable_categories__instant_1ts:mesh = "Mesh2d_face" ;
		colours__mutable_categories__instant_1ts:location = "face" ;
		colours__mutable_categories__instant_1ts:online_operation = "instant" ;
		colours__mutable_categories__instant_1ts:interval_operation = "1 s" ;
		colours__mutable_categories__instant_1ts:interval_write = "1 s" ;
		colours__mutable_categories__instant_1ts:cell_methods = "time: point" ;
		colours__mutable_categories__instant_1ts:coordinates = "time_instant Mesh2d_face_face_y Mesh2d_face_face_x" ;
	double colours__mutable_numbers__instant_1ts(time_counter, mutable_numbers, nMesh2d_face_face) ;
		colours__mutable_numbers__instant_1ts:standard_name = "mutable_numbers" ;
		colours__mutable_numbers__instant_1ts:units = "arbitrary units" ;
		colours__mutable_numbers__instant_1ts:mesh = "Mesh2d_face" ;
		colours__mutable_numbers__instant_1ts:location = "face" ;
		colours__mutable_numbers__instant_1ts:online_operation = "instant" ;
		colours__mutable_numbers__instant_1ts:interval_operation = "1 s" ;
		colours__mutable_numbers__instant_1ts:interval_write = "1 s" ;
		colours__mutable_numbers__instant_1ts:cell_methods = "time: point" ;
		colours__mutable_numbers__instant_1ts:coordinates = "time_instant Mesh2d_face_face_y Mesh2d_face_face_x" ;
	double colours__immutable_both__instant_1ts(time_counter, immutable_numbers, immutable_categories, nMesh2d_face_face) ;
		colours__immutable_both__instant_1ts:standard_name = "immutable_both" ;
		colours__immutable_both__instant_1ts:units = "arbitrary units" ;
		colours__immutable_both__instant_1ts:mesh = "Mesh2d_face" ;
		colours__immutable_both__instant_1ts:location = "face" ;
		colours__immutable_both__instant_1ts:online_operation = "instant" ;
		colours__immutable_both__instant_1ts:interval_operation = "1 s" ;
		colours__immutable_both__instant_1ts:interval_write = "1 s" ;
		colours__immutable_both__instant_1ts:cell_methods = "time: point" ;
		colours__immutable_both__instant_1ts:coordinates = "time_instant Mesh2d_face_face_y Mesh2d_face_face_x" ;

// global attributes:
		:name = "NonSpatialDimensions" ;
		:description = "Created by xios" ;
		:title = "Created by xios" ;
		:Conventions = "UGRID" ;
		:timeStamp = "2021-Aug-20 10:44:46 GMT" ;
		:uuid = "f40b59c8-6f8e-4caa-972c-68bbdba36ba9" ;
data:

 Mesh2d_face_node_x = -45, -15, -15, -45, 15, 15, 45, 45, -45, -15, 15, 45, 
    -45, -15, 15, 45, 75, 75, 105, 105, 135, 135, 75, 105, 135, 75, 105, 135, 
    165, 165, -165, -165, -135, -135, 165, -165, -135, 165, -165, -135, -105, 
    -105, -75, -75, -105, -75, -105, -75, -45, -135, 45, 135, 45, 135, -45, 
    -135 ;

 Mesh2d_face_node_y = 10.72858, 14.51082, 44.00703, 35.26439, 14.51082, 
    44.00703, 10.72858, 35.26439, -10.72858, -14.51082, -14.51082, -10.72858, 
    -35.26439, -44.00703, -44.00703, -35.26439, 14.51082, 44.00703, 14.51082, 
    44.00703, 10.72858, 35.26439, -14.51082, -14.51082, -10.72858, -44.00703, 
    -44.00703, -35.26439, 14.51082, 44.00703, 14.51082, 44.00703, 10.72858, 
    35.26439, -14.51082, -14.51082, -10.72858, -44.00703, -44.00703, 
    -35.26439, 14.51082, 44.00703, 14.51082, 44.00703, -14.51082, -14.51082, 
    -44.00703, -44.00703, 69.24643, 69.24643, 69.24643, 69.24643, -69.24643, 
    -69.24643, -69.24643, -69.24643 ;

 time_instant = 63618879601, 63618879602, 63618879603, 63618879604, 
    63618879605 ;
}
