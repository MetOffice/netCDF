netcdf Fields_grid_nc_C1_T1_201904010000 {
dimensions:
	latitude = 116 ;
	longitude = 122 ;
	nbounds = 2 ;
	string23 = 23 ;
variables:
	float latitude(latitude) ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:axis = "Y" ;
		latitude:valid_min = 48.f ;
		latitude:valid_max = 60.65f ;
		latitude:bounds = "latitude_bounds" ;
	float longitude(longitude) ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:axis = "X" ;
		longitude:valid_min = -11.f ;
		longitude:valid_max = 10.78f ;
		longitude:bounds = "longitude_bounds" ;
	float latitude_bounds(latitude, nbounds) ;
		latitude_bounds:comment = "Bounds" ;
	float longitude_bounds(longitude, nbounds) ;
		longitude_bounds:comment = "Bounds" ;
	int time_0 ;
		time_0:standard_name = "time" ;
		time_0:long_name = "time" ;
		time_0:units = "minutes since 1970-01-01 00:00:00" ;
		time_0:calendar = "gregorian" ;
		time_0:bounds = "time_bnds_0" ;
	int time_bnds_0(nbounds) ;
		time_bnds_0:long_name = "start_and_end_point" ;
	int forecast_reference_time ;
		forecast_reference_time:standard_name = "forecast_reference_time" ;
		forecast_reference_time:long_name = "forecast_reference_time" ;
		forecast_reference_time:units = "minutes since 1970-01-01 00:00:00" ;
		forecast_reference_time:calendar = "gregorian" ;
	int latitude_longitude ;
		latitude_longitude:grid_mapping_name = "latitude_longitude" ;
		latitude_longitude:longitude_of_prime_meridian = 0.f ;
		latitude_longitude:earth_radius = 6371229.f ;
	float height ;
		height:standard_name = "height" ;
		height:comment = "height above ground level" ;
		height:units = "m" ;
		height:long_name = "height above ground level" ;
		height:axis = "Z" ;
		height:positive = "up" ;
		height:reference_datum = "ground level" ;
		height:bounds = "height_bnds" ;
	float height_bnds(nbounds) ;
		height_bnds:long_name = "height above ground level start and end point" ;
	float NO2_CONCENTRATION(latitude, longitude) ;
		NO2_CONCENTRATION:long_name = "NO2_CONCENTRATION" ;
		NO2_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		NO2_CONCENTRATION:field_name = "Unnamed Field Req 1" ;
		NO2_CONCENTRATION:units = "g / m^3" ;
		NO2_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		NO2_CONCENTRATION:quantity = "Concentration" ;
		NO2_CONCENTRATION:species = "NO2" ;
		NO2_CONCENTRATION:species_category = "CHEMISTRY-SPECIES" ;
		NO2_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		NO2_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		NO2_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		NO2_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float O3_CONCENTRATION(latitude, longitude) ;
		O3_CONCENTRATION:long_name = "O3_CONCENTRATION" ;
		O3_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		O3_CONCENTRATION:field_name = "Unnamed Field Req 2" ;
		O3_CONCENTRATION:units = "g / m^3" ;
		O3_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		O3_CONCENTRATION:quantity = "Concentration" ;
		O3_CONCENTRATION:species = "O3" ;
		O3_CONCENTRATION:species_category = "CHEMISTRY-SPECIES" ;
		O3_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		O3_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		O3_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		O3_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float AIT_INS_N_CONCENTRATION(latitude, longitude) ;
		AIT_INS_N_CONCENTRATION:long_name = "AIT_INS_N_CONCENTRATION" ;
		AIT_INS_N_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		AIT_INS_N_CONCENTRATION:field_name = "Unnamed Field Req 3" ;
		AIT_INS_N_CONCENTRATION:units = "1 / m^3" ;
		AIT_INS_N_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		AIT_INS_N_CONCENTRATION:quantity = "Concentration" ;
		AIT_INS_N_CONCENTRATION:species = "Ait_INS_N" ;
		AIT_INS_N_CONCENTRATION:species_category = "CHEMISTRY-SPECIES" ;
		AIT_INS_N_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		AIT_INS_N_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		AIT_INS_N_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		AIT_INS_N_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float AIT_INS_BC_CONCENTRATION(latitude, longitude) ;
		AIT_INS_BC_CONCENTRATION:long_name = "AIT_INS_BC_CONCENTRATION" ;
		AIT_INS_BC_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		AIT_INS_BC_CONCENTRATION:field_name = "Unnamed Field Req 4" ;
		AIT_INS_BC_CONCENTRATION:units = "g / m^3" ;
		AIT_INS_BC_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		AIT_INS_BC_CONCENTRATION:quantity = "Concentration" ;
		AIT_INS_BC_CONCENTRATION:species = "Ait_INS_BC" ;
		AIT_INS_BC_CONCENTRATION:species_category = "CHEMISTRY-SPECIES" ;
		AIT_INS_BC_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		AIT_INS_BC_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		AIT_INS_BC_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		AIT_INS_BC_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float ACC_SOL_SU_CONCENTRATION(latitude, longitude) ;
		ACC_SOL_SU_CONCENTRATION:long_name = "ACC_SOL_SU_CONCENTRATION" ;
		ACC_SOL_SU_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		ACC_SOL_SU_CONCENTRATION:field_name = "Unnamed Field Req 5" ;
		ACC_SOL_SU_CONCENTRATION:units = "g / m^3" ;
		ACC_SOL_SU_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		ACC_SOL_SU_CONCENTRATION:quantity = "Concentration" ;
		ACC_SOL_SU_CONCENTRATION:species = "Acc_SOL_SU" ;
		ACC_SOL_SU_CONCENTRATION:species_category = "CHEMISTRY-SPECIES" ;
		ACC_SOL_SU_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		ACC_SOL_SU_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		ACC_SOL_SU_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		ACC_SOL_SU_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float ACC_SOL_BC_CONCENTRATION(latitude, longitude) ;
		ACC_SOL_BC_CONCENTRATION:long_name = "ACC_SOL_BC_CONCENTRATION" ;
		ACC_SOL_BC_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		ACC_SOL_BC_CONCENTRATION:field_name = "Unnamed Field Req 6" ;
		ACC_SOL_BC_CONCENTRATION:units = "g / m^3" ;
		ACC_SOL_BC_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		ACC_SOL_BC_CONCENTRATION:quantity = "Concentration" ;
		ACC_SOL_BC_CONCENTRATION:species = "Acc_SOL_BC" ;
		ACC_SOL_BC_CONCENTRATION:species_category = "CHEMISTRY-SPECIES" ;
		ACC_SOL_BC_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		ACC_SOL_BC_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		ACC_SOL_BC_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		ACC_SOL_BC_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float ACC_SOL_NH_CONCENTRATION(latitude, longitude) ;
		ACC_SOL_NH_CONCENTRATION:long_name = "ACC_SOL_NH_CONCENTRATION" ;
		ACC_SOL_NH_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		ACC_SOL_NH_CONCENTRATION:field_name = "Unnamed Field Req 7" ;
		ACC_SOL_NH_CONCENTRATION:units = "g / m^3" ;
		ACC_SOL_NH_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		ACC_SOL_NH_CONCENTRATION:quantity = "Concentration" ;
		ACC_SOL_NH_CONCENTRATION:species = "Acc_SOL_NH" ;
		ACC_SOL_NH_CONCENTRATION:species_category = "CHEMISTRY-SPECIES" ;
		ACC_SOL_NH_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		ACC_SOL_NH_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		ACC_SOL_NH_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		ACC_SOL_NH_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float ACC_SOL_NT_CONCENTRATION(latitude, longitude) ;
		ACC_SOL_NT_CONCENTRATION:long_name = "ACC_SOL_NT_CONCENTRATION" ;
		ACC_SOL_NT_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		ACC_SOL_NT_CONCENTRATION:field_name = "Unnamed Field Req 8" ;
		ACC_SOL_NT_CONCENTRATION:units = "g / m^3" ;
		ACC_SOL_NT_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		ACC_SOL_NT_CONCENTRATION:quantity = "Concentration" ;
		ACC_SOL_NT_CONCENTRATION:species = "Acc_SOL_NT" ;
		ACC_SOL_NT_CONCENTRATION:species_category = "CHEMISTRY-SPECIES" ;
		ACC_SOL_NT_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		ACC_SOL_NT_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		ACC_SOL_NT_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		ACC_SOL_NT_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float COR_SOL_SU_CONCENTRATION(latitude, longitude) ;
		COR_SOL_SU_CONCENTRATION:long_name = "COR_SOL_SU_CONCENTRATION" ;
		COR_SOL_SU_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		COR_SOL_SU_CONCENTRATION:field_name = "Unnamed Field Req 9" ;
		COR_SOL_SU_CONCENTRATION:units = "g / m^3" ;
		COR_SOL_SU_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		COR_SOL_SU_CONCENTRATION:quantity = "Concentration" ;
		COR_SOL_SU_CONCENTRATION:species = "Cor_SOL_SU" ;
		COR_SOL_SU_CONCENTRATION:species_category = "CHEMISTRY-SPECIES" ;
		COR_SOL_SU_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		COR_SOL_SU_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		COR_SOL_SU_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		COR_SOL_SU_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float COR_SOL_N_CONCENTRATION(latitude, longitude) ;
		COR_SOL_N_CONCENTRATION:long_name = "COR_SOL_N_CONCENTRATION" ;
		COR_SOL_N_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		COR_SOL_N_CONCENTRATION:field_name = "Unnamed Field Req 10" ;
		COR_SOL_N_CONCENTRATION:units = "1 / m^3" ;
		COR_SOL_N_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		COR_SOL_N_CONCENTRATION:quantity = "Concentration" ;
		COR_SOL_N_CONCENTRATION:species = "Cor_SOL_N" ;
		COR_SOL_N_CONCENTRATION:species_category = "CHEMISTRY-SPECIES" ;
		COR_SOL_N_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		COR_SOL_N_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		COR_SOL_N_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		COR_SOL_N_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float PM10_DRY_CONCENTRATION(latitude, longitude) ;
		PM10_DRY_CONCENTRATION:long_name = "PM10_DRY_CONCENTRATION" ;
		PM10_DRY_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		PM10_DRY_CONCENTRATION:field_name = "Unnamed Field Req 11" ;
		PM10_DRY_CONCENTRATION:units = "g / m^3" ;
		PM10_DRY_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		PM10_DRY_CONCENTRATION:quantity = "Concentration" ;
		PM10_DRY_CONCENTRATION:species = "PM10_dry" ;
		PM10_DRY_CONCENTRATION:species_category = "CHEMISTRY-DIAGN" ;
		PM10_DRY_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		PM10_DRY_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		PM10_DRY_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		PM10_DRY_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float PM2P5_DRY_CONCENTRATION(latitude, longitude) ;
		PM2P5_DRY_CONCENTRATION:long_name = "PM2P5_DRY_CONCENTRATION" ;
		PM2P5_DRY_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		PM2P5_DRY_CONCENTRATION:field_name = "Unnamed Field Req 12" ;
		PM2P5_DRY_CONCENTRATION:units = "g / m^3" ;
		PM2P5_DRY_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		PM2P5_DRY_CONCENTRATION:quantity = "Concentration" ;
		PM2P5_DRY_CONCENTRATION:species = "PM2p5_dry" ;
		PM2P5_DRY_CONCENTRATION:species_category = "CHEMISTRY-DIAGN" ;
		PM2P5_DRY_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		PM2P5_DRY_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		PM2P5_DRY_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		PM2P5_DRY_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float PM10_WET_CONCENTRATION(latitude, longitude) ;
		PM10_WET_CONCENTRATION:long_name = "PM10_WET_CONCENTRATION" ;
		PM10_WET_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		PM10_WET_CONCENTRATION:field_name = "Unnamed Field Req 13" ;
		PM10_WET_CONCENTRATION:units = "g / m^3" ;
		PM10_WET_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		PM10_WET_CONCENTRATION:quantity = "Concentration" ;
		PM10_WET_CONCENTRATION:species = "PM10_wet" ;
		PM10_WET_CONCENTRATION:species_category = "CHEMISTRY-DIAGN" ;
		PM10_WET_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		PM10_WET_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		PM10_WET_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		PM10_WET_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float PM2P5_WET_CONCENTRATION(latitude, longitude) ;
		PM2P5_WET_CONCENTRATION:long_name = "PM2P5_WET_CONCENTRATION" ;
		PM2P5_WET_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		PM2P5_WET_CONCENTRATION:field_name = "Unnamed Field Req 14" ;
		PM2P5_WET_CONCENTRATION:units = "g / m^3" ;
		PM2P5_WET_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		PM2P5_WET_CONCENTRATION:quantity = "Concentration" ;
		PM2P5_WET_CONCENTRATION:species = "PM2p5_wet" ;
		PM2P5_WET_CONCENTRATION:species_category = "CHEMISTRY-DIAGN" ;
		PM2P5_WET_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		PM2P5_WET_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		PM2P5_WET_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		PM2P5_WET_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float PM10_BC_CONCENTRATION(latitude, longitude) ;
		PM10_BC_CONCENTRATION:long_name = "PM10_BC_CONCENTRATION" ;
		PM10_BC_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		PM10_BC_CONCENTRATION:field_name = "Unnamed Field Req 15" ;
		PM10_BC_CONCENTRATION:units = "g / m^3" ;
		PM10_BC_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		PM10_BC_CONCENTRATION:quantity = "Concentration" ;
		PM10_BC_CONCENTRATION:species = "PM10_bc" ;
		PM10_BC_CONCENTRATION:species_category = "CHEMISTRY-DIAGN" ;
		PM10_BC_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		PM10_BC_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		PM10_BC_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		PM10_BC_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float PM2P5_BC_CONCENTRATION(latitude, longitude) ;
		PM2P5_BC_CONCENTRATION:long_name = "PM2P5_BC_CONCENTRATION" ;
		PM2P5_BC_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		PM2P5_BC_CONCENTRATION:field_name = "Unnamed Field Req 16" ;
		PM2P5_BC_CONCENTRATION:units = "g / m^3" ;
		PM2P5_BC_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		PM2P5_BC_CONCENTRATION:quantity = "Concentration" ;
		PM2P5_BC_CONCENTRATION:species = "PM2p5_bc" ;
		PM2P5_BC_CONCENTRATION:species_category = "CHEMISTRY-DIAGN" ;
		PM2P5_BC_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		PM2P5_BC_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		PM2P5_BC_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		PM2P5_BC_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float PM10_OM_CONCENTRATION(latitude, longitude) ;
		PM10_OM_CONCENTRATION:long_name = "PM10_OM_CONCENTRATION" ;
		PM10_OM_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		PM10_OM_CONCENTRATION:field_name = "Unnamed Field Req 17" ;
		PM10_OM_CONCENTRATION:units = "g / m^3" ;
		PM10_OM_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		PM10_OM_CONCENTRATION:quantity = "Concentration" ;
		PM10_OM_CONCENTRATION:species = "PM10_om" ;
		PM10_OM_CONCENTRATION:species_category = "CHEMISTRY-DIAGN" ;
		PM10_OM_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		PM10_OM_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		PM10_OM_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		PM10_OM_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float PM2P5_OM_CONCENTRATION(latitude, longitude) ;
		PM2P5_OM_CONCENTRATION:long_name = "PM2P5_OM_CONCENTRATION" ;
		PM2P5_OM_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		PM2P5_OM_CONCENTRATION:field_name = "Unnamed Field Req 18" ;
		PM2P5_OM_CONCENTRATION:units = "g / m^3" ;
		PM2P5_OM_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		PM2P5_OM_CONCENTRATION:quantity = "Concentration" ;
		PM2P5_OM_CONCENTRATION:species = "PM2p5_om" ;
		PM2P5_OM_CONCENTRATION:species_category = "CHEMISTRY-DIAGN" ;
		PM2P5_OM_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		PM2P5_OM_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		PM2P5_OM_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		PM2P5_OM_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float PM10_H2SO4_CONCENTRATION(latitude, longitude) ;
		PM10_H2SO4_CONCENTRATION:long_name = "PM10_H2SO4_CONCENTRATION" ;
		PM10_H2SO4_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		PM10_H2SO4_CONCENTRATION:field_name = "Unnamed Field Req 19" ;
		PM10_H2SO4_CONCENTRATION:units = "g / m^3" ;
		PM10_H2SO4_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		PM10_H2SO4_CONCENTRATION:quantity = "Concentration" ;
		PM10_H2SO4_CONCENTRATION:species = "PM10_h2so4" ;
		PM10_H2SO4_CONCENTRATION:species_category = "CHEMISTRY-DIAGN" ;
		PM10_H2SO4_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		PM10_H2SO4_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		PM10_H2SO4_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		PM10_H2SO4_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float PM2P5_H2SO4_CONCENTRATION(latitude, longitude) ;
		PM2P5_H2SO4_CONCENTRATION:long_name = "PM2P5_H2SO4_CONCENTRATION" ;
		PM2P5_H2SO4_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		PM2P5_H2SO4_CONCENTRATION:field_name = "Unnamed Field Req 20" ;
		PM2P5_H2SO4_CONCENTRATION:units = "g / m^3" ;
		PM2P5_H2SO4_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		PM2P5_H2SO4_CONCENTRATION:quantity = "Concentration" ;
		PM2P5_H2SO4_CONCENTRATION:species = "PM2p5_h2so4" ;
		PM2P5_H2SO4_CONCENTRATION:species_category = "CHEMISTRY-DIAGN" ;
		PM2P5_H2SO4_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		PM2P5_H2SO4_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		PM2P5_H2SO4_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		PM2P5_H2SO4_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float PM10_SS_CONCENTRATION(latitude, longitude) ;
		PM10_SS_CONCENTRATION:long_name = "PM10_SS_CONCENTRATION" ;
		PM10_SS_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		PM10_SS_CONCENTRATION:field_name = "Unnamed Field Req 21" ;
		PM10_SS_CONCENTRATION:units = "g / m^3" ;
		PM10_SS_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		PM10_SS_CONCENTRATION:quantity = "Concentration" ;
		PM10_SS_CONCENTRATION:species = "PM10_ss" ;
		PM10_SS_CONCENTRATION:species_category = "CHEMISTRY-DIAGN" ;
		PM10_SS_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		PM10_SS_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		PM10_SS_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		PM10_SS_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float PM2P5_SS_CONCENTRATION(latitude, longitude) ;
		PM2P5_SS_CONCENTRATION:long_name = "PM2P5_SS_CONCENTRATION" ;
		PM2P5_SS_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		PM2P5_SS_CONCENTRATION:field_name = "Unnamed Field Req 22" ;
		PM2P5_SS_CONCENTRATION:units = "g / m^3" ;
		PM2P5_SS_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		PM2P5_SS_CONCENTRATION:quantity = "Concentration" ;
		PM2P5_SS_CONCENTRATION:species = "PM2p5_ss" ;
		PM2P5_SS_CONCENTRATION:species_category = "CHEMISTRY-DIAGN" ;
		PM2P5_SS_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		PM2P5_SS_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		PM2P5_SS_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		PM2P5_SS_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float PM10_NH4_CONCENTRATION(latitude, longitude) ;
		PM10_NH4_CONCENTRATION:long_name = "PM10_NH4_CONCENTRATION" ;
		PM10_NH4_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		PM10_NH4_CONCENTRATION:field_name = "Unnamed Field Req 23" ;
		PM10_NH4_CONCENTRATION:units = "g / m^3" ;
		PM10_NH4_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		PM10_NH4_CONCENTRATION:quantity = "Concentration" ;
		PM10_NH4_CONCENTRATION:species = "PM10_nh4" ;
		PM10_NH4_CONCENTRATION:species_category = "CHEMISTRY-DIAGN" ;
		PM10_NH4_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		PM10_NH4_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		PM10_NH4_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		PM10_NH4_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float PM2P5_NH4_CONCENTRATION(latitude, longitude) ;
		PM2P5_NH4_CONCENTRATION:long_name = "PM2P5_NH4_CONCENTRATION" ;
		PM2P5_NH4_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		PM2P5_NH4_CONCENTRATION:field_name = "Unnamed Field Req 24" ;
		PM2P5_NH4_CONCENTRATION:units = "g / m^3" ;
		PM2P5_NH4_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		PM2P5_NH4_CONCENTRATION:quantity = "Concentration" ;
		PM2P5_NH4_CONCENTRATION:species = "PM2p5_nh4" ;
		PM2P5_NH4_CONCENTRATION:species_category = "CHEMISTRY-DIAGN" ;
		PM2P5_NH4_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		PM2P5_NH4_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		PM2P5_NH4_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		PM2P5_NH4_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float PM10_NO3_CONCENTRATION(latitude, longitude) ;
		PM10_NO3_CONCENTRATION:long_name = "PM10_NO3_CONCENTRATION" ;
		PM10_NO3_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		PM10_NO3_CONCENTRATION:field_name = "Unnamed Field Req 25" ;
		PM10_NO3_CONCENTRATION:units = "g / m^3" ;
		PM10_NO3_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		PM10_NO3_CONCENTRATION:quantity = "Concentration" ;
		PM10_NO3_CONCENTRATION:species = "PM10_no3" ;
		PM10_NO3_CONCENTRATION:species_category = "CHEMISTRY-DIAGN" ;
		PM10_NO3_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		PM10_NO3_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		PM10_NO3_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		PM10_NO3_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float PM2P5_NO3_CONCENTRATION(latitude, longitude) ;
		PM2P5_NO3_CONCENTRATION:long_name = "PM2P5_NO3_CONCENTRATION" ;
		PM2P5_NO3_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		PM2P5_NO3_CONCENTRATION:field_name = "Unnamed Field Req 26" ;
		PM2P5_NO3_CONCENTRATION:units = "g / m^3" ;
		PM2P5_NO3_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		PM2P5_NO3_CONCENTRATION:quantity = "Concentration" ;
		PM2P5_NO3_CONCENTRATION:species = "PM2p5_no3" ;
		PM2P5_NO3_CONCENTRATION:species_category = "CHEMISTRY-DIAGN" ;
		PM2P5_NO3_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		PM2P5_NO3_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		PM2P5_NO3_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		PM2P5_NO3_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float PM10_NN_CONCENTRATION(latitude, longitude) ;
		PM10_NN_CONCENTRATION:long_name = "PM10_NN_CONCENTRATION" ;
		PM10_NN_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		PM10_NN_CONCENTRATION:field_name = "Unnamed Field Req 27" ;
		PM10_NN_CONCENTRATION:units = "g / m^3" ;
		PM10_NN_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		PM10_NN_CONCENTRATION:quantity = "Concentration" ;
		PM10_NN_CONCENTRATION:species = "PM10_nn" ;
		PM10_NN_CONCENTRATION:species_category = "CHEMISTRY-DIAGN" ;
		PM10_NN_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		PM10_NN_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		PM10_NN_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		PM10_NN_CONCENTRATION:cell_methods = "time: mean height: mean" ;
	float PM2P5_NN_CONCENTRATION(latitude, longitude) ;
		PM2P5_NN_CONCENTRATION:long_name = "PM2P5_NN_CONCENTRATION" ;
		PM2P5_NN_CONCENTRATION:grid_mapping = "latitude_longitude" ;
		PM2P5_NN_CONCENTRATION:field_name = "Unnamed Field Req 28" ;
		PM2P5_NN_CONCENTRATION:units = "g / m^3" ;
		PM2P5_NN_CONCENTRATION:coordinates = "time_0 forecast_reference_time height" ;
		PM2P5_NN_CONCENTRATION:quantity = "Concentration" ;
		PM2P5_NN_CONCENTRATION:species = "PM2p5_nn" ;
		PM2P5_NN_CONCENTRATION:species_category = "CHEMISTRY-DIAGN" ;
		PM2P5_NN_CONCENTRATION:time_av_int_info = "1hr 0min average" ;
		PM2P5_NN_CONCENTRATION:vertical_av_int_info = "Finite Z-average" ;
		PM2P5_NN_CONCENTRATION:horizontal_av_int_info = "No horizontal averaging" ;
		PM2P5_NN_CONCENTRATION:cell_methods = "time: mean height: mean" ;

// global attributes:
		:title = "Scientific - Eulerian AQ UKCA RAQ MODE 10" ;
		:Conventions = "CF-1.8" ;
		:history = "NAME 13/11/2025 15:44:09.178 UTC" ;
		:source = "Met Office NAME model" ;
		:institution = "NA" ;
		:reference = "https://doi.org/10.1007/978-0-387-68854-1_62" ;
		:comment = "none" ;
		:name_version = "NAME III (development version 8.7+)" ;
		:run_time = "13/11/2025 15:44:09.178 UTC" ;
		:run_duration = "358577day 0hr 0min" ;
		:met_data = "NWP Flow.Regional" ;
		:name_netcdf_out_vers = "0.1" ;
		:start_of_release = "-infinity" ;
		:end_of_release = "infinity" ;
		:source_strength = "Multiple Sources" ;
		:release_location = "Multiple Sources" ;
		:release_height = "Multiple Sources" ;
}
