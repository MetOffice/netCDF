netcdf \20210315T0700Z-PT0001H00M-precip_rate {
dimensions:
	threshold = 12 ;
	latitude = 960 ;
	longitude = 1280 ;
	bnds = 2 ;
variables:
	float probability_of_lwe_precipitation_rate_above_threshold(threshold, latitude, longitude) ;
		probability_of_lwe_precipitation_rate_above_threshold:long_name = "probability_of_lwe_precipitation_rate_above_threshold" ;
		probability_of_lwe_precipitation_rate_above_threshold:units = "1" ;
		probability_of_lwe_precipitation_rate_above_threshold:grid_mapping = "latitude_longitude" ;
		probability_of_lwe_precipitation_rate_above_threshold:coordinates = "blend_time forecast_period forecast_reference_time time" ;
	int latitude_longitude ;
		latitude_longitude:grid_mapping_name = "latitude_longitude" ;
		latitude_longitude:longitude_of_prime_meridian = 0. ;
		latitude_longitude:earth_radius = 6371229. ;
	float threshold(threshold) ;
		threshold:units = "m s-1" ;
		threshold:standard_name = "lwe_precipitation_rate" ;
		threshold:spp__relative_to_threshold = "greater_than" ;
	float latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:bounds = "latitude_bnds" ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
	float latitude_bnds(latitude, bnds) ;
	float longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:bounds = "longitude_bnds" ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;
	float longitude_bnds(longitude, bnds) ;
	int64 blend_time ;
		blend_time:units = "seconds since 1970-01-01 00:00:00" ;
		blend_time:long_name = "blend_time" ;
		blend_time:calendar = "gregorian" ;
	int forecast_period ;
		forecast_period:units = "seconds" ;
		forecast_period:standard_name = "forecast_period" ;
		forecast_period:deprecation_message = "forecast_period will be removed in future and should not be used" ;
	int64 forecast_reference_time ;
		forecast_reference_time:units = "seconds since 1970-01-01 00:00:00" ;
		forecast_reference_time:standard_name = "forecast_reference_time" ;
		forecast_reference_time:calendar = "gregorian" ;
		forecast_reference_time:deprecation_message = "forecast_reference_time will be removed in future and should not be used" ;
	int64 time ;
		time:units = "seconds since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "gregorian" ;

// global attributes:
		:institution = "Met Office" ;
		:mosg__model_configuration = "gl_ens" ;
		:source = "Met Office Unified Model" ;
		:title = "Post-Processed MOGREPS-G Model Forecast on Global 20 km Standard Grid" ;
		:Conventions = "CF-1.5" ;
data:

 threshold = 0, 8.333333e-09, 2.777778e-08, 6.944445e-08, 1.388889e-07, 
    2.777778e-07, 5.555556e-07, 1.111111e-06, 2.222222e-06, 4.444445e-06, 
    8.888889e-06, 1.777778e-05 ;

 time = 1615791600 ;
}
